module ADDER (
\data1_in[0], 
\data1_in[10], 
\data1_in[11], 
\data1_in[12], 
\data1_in[13], 
\data1_in[14], 
\data1_in[15], 
\data1_in[16], 
\data1_in[17], 
\data1_in[18], 
\data1_in[19], 
\data1_in[1], 
\data1_in[20], 
\data1_in[21], 
\data1_in[22], 
\data1_in[23], 
\data1_in[24], 
\data1_in[25], 
\data1_in[26], 
\data1_in[27], 
\data1_in[28], 
\data1_in[29], 
\data1_in[2], 
\data1_in[30], 
\data1_in[31], 
\data1_in[3], 
\data1_in[4], 
\data1_in[5], 
\data1_in[6], 
\data1_in[7], 
\data1_in[8], 
\data1_in[9], 
\data2_in[0], 
\data2_in[10], 
\data2_in[11], 
\data2_in[12], 
\data2_in[13], 
\data2_in[14], 
\data2_in[15], 
\data2_in[16], 
\data2_in[17], 
\data2_in[18], 
\data2_in[19], 
\data2_in[1], 
\data2_in[20], 
\data2_in[21], 
\data2_in[22], 
\data2_in[23], 
\data2_in[24], 
\data2_in[25], 
\data2_in[26], 
\data2_in[27], 
\data2_in[28], 
\data2_in[29], 
\data2_in[2], 
\data2_in[30], 
\data2_in[31], 
\data2_in[3], 
\data2_in[4], 
\data2_in[5], 
\data2_in[6], 
\data2_in[7], 
\data2_in[8], 
\data2_in[9],
\data_o[0], 
\data_o[10], 
\data_o[11], 
\data_o[12], 
\data_o[13], 
\data_o[14], 
\data_o[15], 
\data_o[16], 
\data_o[17], 
\data_o[18], 
\data_o[19], 
\data_o[1], 
\data_o[20], 
\data_o[21], 
\data_o[22], 
\data_o[23], 
\data_o[24], 
\data_o[25], 
\data_o[26], 
\data_o[27], 
\data_o[28], 
\data_o[29], 
\data_o[2], 
\data_o[30], 
\data_o[31], 
\data_o[3], 
\data_o[4], 
\data_o[5], 
\data_o[6], 
\data_o[7], 
\data_o[8], 
\data_o[9]
);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  input \data1_in[0];
  input \data1_in[10];
  input \data1_in[11];
  input \data1_in[12];
  input \data1_in[13];
  input \data1_in[14];
  input \data1_in[15];
  input \data1_in[16];
  input \data1_in[17];
  input \data1_in[18];
  input \data1_in[19];
  input \data1_in[1];
  input \data1_in[20];
  input \data1_in[21];
  input \data1_in[22];
  input \data1_in[23];
  input \data1_in[24];
  input \data1_in[25];
  input \data1_in[26];
  input \data1_in[27];
  input \data1_in[28];
  input \data1_in[29];
  input \data1_in[2];
  input \data1_in[30];
  input \data1_in[31];
  input \data1_in[3];
  input \data1_in[4];
  input \data1_in[5];
  input \data1_in[6];
  input \data1_in[7];
  input \data1_in[8];
  input \data1_in[9];
  input \data2_in[0];
  input \data2_in[10];
  input \data2_in[11];
  input \data2_in[12];
  input \data2_in[13];
  input \data2_in[14];
  input \data2_in[15];
  input \data2_in[16];
  input \data2_in[17];
  input \data2_in[18];
  input \data2_in[19];
  input \data2_in[1];
  input \data2_in[20];
  input \data2_in[21];
  input \data2_in[22];
  input \data2_in[23];
  input \data2_in[24];
  input \data2_in[25];
  input \data2_in[26];
  input \data2_in[27];
  input \data2_in[28];
  input \data2_in[29];
  input \data2_in[2];
  input \data2_in[30];
  input \data2_in[31];
  input \data2_in[3];
  input \data2_in[4];
  input \data2_in[5];
  input \data2_in[6];
  input \data2_in[7];
  input \data2_in[8];
  input \data2_in[9];
  output \data_o[0];
  output \data_o[10];
  output \data_o[11];
  output \data_o[12];
  output \data_o[13];
  output \data_o[14];
  output \data_o[15];
  output \data_o[16];
  output \data_o[17];
  output \data_o[18];
  output \data_o[19];
  output \data_o[1];
  output \data_o[20];
  output \data_o[21];
  output \data_o[22];
  output \data_o[23];
  output \data_o[24];
  output \data_o[25];
  output \data_o[26];
  output \data_o[27];
  output \data_o[28];
  output \data_o[29];
  output \data_o[2];
  output \data_o[30];
  output \data_o[31];
  output \data_o[3];
  output \data_o[4];
  output \data_o[5];
  output \data_o[6];
  output \data_o[7];
  output \data_o[8];
  output \data_o[9];
  NAND _137_ (
    .A(\data2_in[14] ),
    .B(\data1_in[14] ),
    .Y(_134_)
  );
  XOR _138_ (
    .A(\data2_in[14] ),
    .B(\data1_in[14] ),
    .Y(_135_)
  );
  OR _139_ (
    .A(\data2_in[13] ),
    .B(\data1_in[13] ),
    .Y(_136_)
  );
  NAND _140_ (
    .A(\data2_in[12] ),
    .B(\data1_in[12] ),
    .Y(_000_)
  );
  XOR _141_ (
    .A(\data2_in[12] ),
    .B(\data1_in[12] ),
    .Y(_001_)
  );
  NAND _142_ (
    .A(\data2_in[11] ),
    .B(\data1_in[11] ),
    .Y(_002_)
  );
  OR _143_ (
    .A(\data2_in[11] ),
    .B(\data1_in[11] ),
    .Y(_003_)
  );
  NAND _144_ (
    .A(\data2_in[10] ),
    .B(\data1_in[10] ),
    .Y(_004_)
  );
  XOR _145_ (
    .A(\data2_in[10] ),
    .B(\data1_in[10] ),
    .Y(_005_)
  );
  OR _146_ (
    .A(\data2_in[9] ),
    .B(\data1_in[9] ),
    .Y(_006_)
  );
  NAND _147_ (
    .A(\data2_in[9] ),
    .B(\data1_in[9] ),
    .Y(_007_)
  );
  NAND _148_ (
    .A(\data2_in[8] ),
    .B(\data1_in[8] ),
    .Y(_008_)
  );
  XOR _149_ (
    .A(\data2_in[8] ),
    .B(\data1_in[8] ),
    .Y(_009_)
  );
  NAND _150_ (
    .A(\data2_in[7] ),
    .B(\data1_in[7] ),
    .Y(_010_)
  );
  OR _151_ (
    .A(\data2_in[7] ),
    .B(\data1_in[7] ),
    .Y(_011_)
  );
  NAND _152_ (
    .A(\data2_in[6] ),
    .B(\data1_in[6] ),
    .Y(_012_)
  );
  XOR _153_ (
    .A(\data2_in[6] ),
    .B(\data1_in[6] ),
    .Y(_013_)
  );
  NAND _154_ (
    .A(\data2_in[5] ),
    .B(\data1_in[5] ),
    .Y(_014_)
  );
  OR _155_ (
    .A(\data2_in[5] ),
    .B(\data1_in[5] ),
    .Y(_015_)
  );
  NAND _156_ (
    .A(\data2_in[4] ),
    .B(\data1_in[4] ),
    .Y(_016_)
  );
  XOR _157_ (
    .A(\data2_in[4] ),
    .B(\data1_in[4] ),
    .Y(_017_)
  );
  NAND _158_ (
    .A(\data2_in[3] ),
    .B(\data1_in[3] ),
    .Y(_018_)
  );
  OR _159_ (
    .A(\data2_in[3] ),
    .B(\data1_in[3] ),
    .Y(_019_)
  );
  NAND _160_ (
    .A(\data2_in[2] ),
    .B(\data1_in[2] ),
    .Y(_020_)
  );
  NAND _161_ (
    .A(\data2_in[1] ),
    .B(\data1_in[1] ),
    .Y(_021_)
  );
  AND _162_ (
    .A(\data2_in[0] ),
    .B(\data1_in[0] ),
    .Y(_022_)
  );
  XOR _163_ (
    .A(\data2_in[1] ),
    .B(\data1_in[1] ),
    .Y(_023_)
  );
  NAND _164_ (
    .A(_022_),
    .B(_023_),
    .Y(_024_)
  );
  NAND _165_ (
    .A(_021_),
    .B(_024_),
    .Y(_025_)
  );
  XOR _166_ (
    .A(\data2_in[2] ),
    .B(\data1_in[2] ),
    .Y(_026_)
  );
  NAND _167_ (
    .A(_025_),
    .B(_026_),
    .Y(_027_)
  );
  NAND _168_ (
    .A(_020_),
    .B(_027_),
    .Y(_028_)
  );
  NAND _169_ (
    .A(_019_),
    .B(_028_),
    .Y(_029_)
  );
  NAND _170_ (
    .A(_018_),
    .B(_029_),
    .Y(_030_)
  );
  NAND _171_ (
    .A(_017_),
    .B(_030_),
    .Y(_031_)
  );
  NAND _172_ (
    .A(_016_),
    .B(_031_),
    .Y(_032_)
  );
  NAND _173_ (
    .A(_015_),
    .B(_032_),
    .Y(_033_)
  );
  NAND _174_ (
    .A(_014_),
    .B(_033_),
    .Y(_034_)
  );
  NAND _175_ (
    .A(_013_),
    .B(_034_),
    .Y(_035_)
  );
  NAND _176_ (
    .A(_012_),
    .B(_035_),
    .Y(_036_)
  );
  NAND _177_ (
    .A(_011_),
    .B(_036_),
    .Y(_037_)
  );
  NAND _178_ (
    .A(_010_),
    .B(_037_),
    .Y(_038_)
  );
  NAND _179_ (
    .A(_009_),
    .B(_038_),
    .Y(_039_)
  );
  AND _180_ (
    .A(_008_),
    .B(_039_),
    .Y(_040_)
  );
  NAND _181_ (
    .A(_007_),
    .B(_040_),
    .Y(_041_)
  );
  AND _182_ (
    .A(_006_),
    .B(_041_),
    .Y(_042_)
  );
  NAND _183_ (
    .A(_005_),
    .B(_042_),
    .Y(_043_)
  );
  NAND _184_ (
    .A(_004_),
    .B(_043_),
    .Y(_044_)
  );
  NAND _185_ (
    .A(_003_),
    .B(_044_),
    .Y(_045_)
  );
  NAND _186_ (
    .A(_002_),
    .B(_045_),
    .Y(_046_)
  );
  NAND _187_ (
    .A(_001_),
    .B(_046_),
    .Y(_047_)
  );
  NAND _188_ (
    .A(\data2_in[13] ),
    .B(\data1_in[13] ),
    .Y(_048_)
  );
  AND _189_ (
    .A(_000_),
    .B(_048_),
    .Y(_049_)
  );
  NAND _190_ (
    .A(_047_),
    .B(_049_),
    .Y(_050_)
  );
  AND _191_ (
    .A(_136_),
    .B(_048_),
    .Y(_051_)
  );
  AND _192_ (
    .A(_136_),
    .B(_050_),
    .Y(_052_)
  );
  NAND _193_ (
    .A(_135_),
    .B(_052_),
    .Y(_053_)
  );
  XOR _194_ (
    .A(_135_),
    .B(_052_),
    .Y(\data_o[14] )
  );
  NAND _195_ (
    .A(_134_),
    .B(_053_),
    .Y(_054_)
  );
  NAND _196_ (
    .A(\data2_in[15] ),
    .B(\data1_in[15] ),
    .Y(_055_)
  );
  OR _197_ (
    .A(\data2_in[15] ),
    .B(\data1_in[15] ),
    .Y(_056_)
  );
  AND _198_ (
    .A(_055_),
    .B(_056_),
    .Y(_057_)
  );
  XOR _199_ (
    .A(_054_),
    .B(_057_),
    .Y(\data_o[15] )
  );
  NAND _200_ (
    .A(\data2_in[16] ),
    .B(\data1_in[16] ),
    .Y(_058_)
  );
  XOR _201_ (
    .A(\data2_in[16] ),
    .B(\data1_in[16] ),
    .Y(_059_)
  );
  AND _202_ (
    .A(_134_),
    .B(_055_),
    .Y(_060_)
  );
  NAND _203_ (
    .A(_053_),
    .B(_060_),
    .Y(_061_)
  );
  AND _204_ (
    .A(_056_),
    .B(_061_),
    .Y(_062_)
  );
  NAND _205_ (
    .A(_059_),
    .B(_062_),
    .Y(_063_)
  );
  XOR _206_ (
    .A(_059_),
    .B(_062_),
    .Y(\data_o[16] )
  );
  NAND _207_ (
    .A(_058_),
    .B(_063_),
    .Y(_064_)
  );
  NAND _208_ (
    .A(\data2_in[17] ),
    .B(\data1_in[17] ),
    .Y(_065_)
  );
  OR _209_ (
    .A(\data2_in[17] ),
    .B(\data1_in[17] ),
    .Y(_066_)
  );
  AND _210_ (
    .A(_065_),
    .B(_066_),
    .Y(_067_)
  );
  XOR _211_ (
    .A(_064_),
    .B(_067_),
    .Y(\data_o[17] )
  );
  NAND _212_ (
    .A(\data2_in[18] ),
    .B(\data1_in[18] ),
    .Y(_068_)
  );
  XOR _213_ (
    .A(\data2_in[18] ),
    .B(\data1_in[18] ),
    .Y(_069_)
  );
  AND _214_ (
    .A(_058_),
    .B(_065_),
    .Y(_070_)
  );
  NAND _215_ (
    .A(_063_),
    .B(_070_),
    .Y(_071_)
  );
  AND _216_ (
    .A(_066_),
    .B(_071_),
    .Y(_072_)
  );
  NAND _217_ (
    .A(_069_),
    .B(_072_),
    .Y(_073_)
  );
  XOR _218_ (
    .A(_069_),
    .B(_072_),
    .Y(\data_o[18] )
  );
  NAND _219_ (
    .A(_068_),
    .B(_073_),
    .Y(_074_)
  );
  NAND _220_ (
    .A(\data2_in[19] ),
    .B(\data1_in[19] ),
    .Y(_075_)
  );
  OR _221_ (
    .A(\data2_in[19] ),
    .B(\data1_in[19] ),
    .Y(_076_)
  );
  AND _222_ (
    .A(_075_),
    .B(_076_),
    .Y(_077_)
  );
  XOR _223_ (
    .A(_074_),
    .B(_077_),
    .Y(\data_o[19] )
  );
  NAND _224_ (
    .A(\data2_in[20] ),
    .B(\data1_in[20] ),
    .Y(_078_)
  );
  XOR _225_ (
    .A(\data2_in[20] ),
    .B(\data1_in[20] ),
    .Y(_079_)
  );
  NAND _226_ (
    .A(_074_),
    .B(_076_),
    .Y(_080_)
  );
  NAND _227_ (
    .A(_075_),
    .B(_080_),
    .Y(_081_)
  );
  NAND _228_ (
    .A(_079_),
    .B(_081_),
    .Y(_082_)
  );
  XOR _229_ (
    .A(_079_),
    .B(_081_),
    .Y(\data_o[20] )
  );
  NAND _230_ (
    .A(_078_),
    .B(_082_),
    .Y(_083_)
  );
  NAND _231_ (
    .A(\data2_in[21] ),
    .B(\data1_in[21] ),
    .Y(_084_)
  );
  OR _232_ (
    .A(\data2_in[21] ),
    .B(\data1_in[21] ),
    .Y(_085_)
  );
  AND _233_ (
    .A(_084_),
    .B(_085_),
    .Y(_086_)
  );
  XOR _234_ (
    .A(_083_),
    .B(_086_),
    .Y(\data_o[21] )
  );
  NAND _235_ (
    .A(\data2_in[22] ),
    .B(\data1_in[22] ),
    .Y(_087_)
  );
  XOR _236_ (
    .A(\data2_in[22] ),
    .B(\data1_in[22] ),
    .Y(_088_)
  );
  NAND _237_ (
    .A(_083_),
    .B(_085_),
    .Y(_089_)
  );
  NAND _238_ (
    .A(_084_),
    .B(_089_),
    .Y(_090_)
  );
  NAND _239_ (
    .A(_088_),
    .B(_090_),
    .Y(_091_)
  );
  XOR _240_ (
    .A(_088_),
    .B(_090_),
    .Y(\data_o[22] )
  );
  NAND _241_ (
    .A(_087_),
    .B(_091_),
    .Y(_092_)
  );
  NAND _242_ (
    .A(\data2_in[23] ),
    .B(\data1_in[23] ),
    .Y(_093_)
  );
  OR _243_ (
    .A(\data2_in[23] ),
    .B(\data1_in[23] ),
    .Y(_094_)
  );
  AND _244_ (
    .A(_093_),
    .B(_094_),
    .Y(_095_)
  );
  XOR _245_ (
    .A(_092_),
    .B(_095_),
    .Y(\data_o[23] )
  );
  NAND _246_ (
    .A(\data2_in[24] ),
    .B(\data1_in[24] ),
    .Y(_096_)
  );
  XOR _247_ (
    .A(\data2_in[24] ),
    .B(\data1_in[24] ),
    .Y(_097_)
  );
  NAND _248_ (
    .A(_092_),
    .B(_094_),
    .Y(_098_)
  );
  NAND _249_ (
    .A(_093_),
    .B(_098_),
    .Y(_099_)
  );
  NAND _250_ (
    .A(_097_),
    .B(_099_),
    .Y(_100_)
  );
  XOR _251_ (
    .A(_097_),
    .B(_099_),
    .Y(\data_o[24] )
  );
  NAND _252_ (
    .A(_096_),
    .B(_100_),
    .Y(_101_)
  );
  NAND _253_ (
    .A(\data2_in[25] ),
    .B(\data1_in[25] ),
    .Y(_102_)
  );
  XOR _254_ (
    .A(\data2_in[25] ),
    .B(\data1_in[25] ),
    .Y(_103_)
  );
  NAND _255_ (
    .A(_101_),
    .B(_103_),
    .Y(_104_)
  );
  XOR _256_ (
    .A(_101_),
    .B(_103_),
    .Y(\data_o[25] )
  );
  NAND _257_ (
    .A(_102_),
    .B(_104_),
    .Y(_105_)
  );
  NAND _258_ (
    .A(\data2_in[26] ),
    .B(\data1_in[26] ),
    .Y(_106_)
  );
  XOR _259_ (
    .A(\data2_in[26] ),
    .B(\data1_in[26] ),
    .Y(_107_)
  );
  NAND _260_ (
    .A(_105_),
    .B(_107_),
    .Y(_108_)
  );
  XOR _261_ (
    .A(_105_),
    .B(_107_),
    .Y(\data_o[26] )
  );
  NAND _262_ (
    .A(_106_),
    .B(_108_),
    .Y(_109_)
  );
  NAND _263_ (
    .A(\data2_in[27] ),
    .B(\data1_in[27] ),
    .Y(_110_)
  );
  OR _264_ (
    .A(\data2_in[27] ),
    .B(\data1_in[27] ),
    .Y(_111_)
  );
  AND _265_ (
    .A(_110_),
    .B(_111_),
    .Y(_112_)
  );
  XOR _266_ (
    .A(_109_),
    .B(_112_),
    .Y(\data_o[27] )
  );
  NAND _267_ (
    .A(\data2_in[28] ),
    .B(\data1_in[28] ),
    .Y(_113_)
  );
  XOR _268_ (
    .A(\data2_in[28] ),
    .B(\data1_in[28] ),
    .Y(_114_)
  );
  NAND _269_ (
    .A(_109_),
    .B(_111_),
    .Y(_115_)
  );
  NAND _270_ (
    .A(_110_),
    .B(_115_),
    .Y(_116_)
  );
  NAND _271_ (
    .A(_114_),
    .B(_116_),
    .Y(_117_)
  );
  XOR _272_ (
    .A(_114_),
    .B(_116_),
    .Y(\data_o[28] )
  );
  NAND _273_ (
    .A(_113_),
    .B(_117_),
    .Y(_118_)
  );
  NAND _274_ (
    .A(\data2_in[29] ),
    .B(\data1_in[29] ),
    .Y(_119_)
  );
  XOR _275_ (
    .A(\data2_in[29] ),
    .B(\data1_in[29] ),
    .Y(_120_)
  );
  NAND _276_ (
    .A(_118_),
    .B(_120_),
    .Y(_121_)
  );
  XOR _277_ (
    .A(_118_),
    .B(_120_),
    .Y(\data_o[29] )
  );
  NAND _278_ (
    .A(_119_),
    .B(_121_),
    .Y(_122_)
  );
  NAND _279_ (
    .A(\data2_in[30] ),
    .B(\data1_in[30] ),
    .Y(_123_)
  );
  XOR _280_ (
    .A(\data2_in[30] ),
    .B(\data1_in[30] ),
    .Y(_124_)
  );
  NAND _281_ (
    .A(_122_),
    .B(_124_),
    .Y(_125_)
  );
  XOR _282_ (
    .A(_122_),
    .B(_124_),
    .Y(\data_o[30] )
  );
  NAND _283_ (
    .A(_123_),
    .B(_125_),
    .Y(_126_)
  );
  XOR _284_ (
    .A(\data2_in[31] ),
    .B(\data1_in[31] ),
    .Y(_127_)
  );
  XOR _285_ (
    .A(_126_),
    .B(_127_),
    .Y(\data_o[31] )
  );
  XOR _286_ (
    .A(\data2_in[0] ),
    .B(\data1_in[0] ),
    .Y(\data_o[0] )
  );
  XOR _287_ (
    .A(_022_),
    .B(_023_),
    .Y(\data_o[1] )
  );
  XOR _288_ (
    .A(_025_),
    .B(_026_),
    .Y(\data_o[2] )
  );
  AND _289_ (
    .A(_018_),
    .B(_019_),
    .Y(_128_)
  );
  XOR _290_ (
    .A(_028_),
    .B(_128_),
    .Y(\data_o[3] )
  );
  XOR _291_ (
    .A(_017_),
    .B(_030_),
    .Y(\data_o[4] )
  );
  AND _292_ (
    .A(_014_),
    .B(_015_),
    .Y(_129_)
  );
  XOR _293_ (
    .A(_032_),
    .B(_129_),
    .Y(\data_o[5] )
  );
  XOR _294_ (
    .A(_013_),
    .B(_034_),
    .Y(\data_o[6] )
  );
  AND _295_ (
    .A(_010_),
    .B(_011_),
    .Y(_130_)
  );
  XOR _296_ (
    .A(_036_),
    .B(_130_),
    .Y(\data_o[7] )
  );
  XOR _297_ (
    .A(_009_),
    .B(_038_),
    .Y(\data_o[8] )
  );
  NAND _298_ (
    .A(_006_),
    .B(_007_),
    .Y(_131_)
  );
  XOR _299_ (
    .A(_040_),
    .B(_131_),
    .Y(\data_o[9] )
  );
  XOR _300_ (
    .A(_005_),
    .B(_042_),
    .Y(\data_o[10] )
  );
  AND _301_ (
    .A(_002_),
    .B(_003_),
    .Y(_132_)
  );
  XOR _302_ (
    .A(_044_),
    .B(_132_),
    .Y(\data_o[11] )
  );
  XOR _303_ (
    .A(_001_),
    .B(_046_),
    .Y(\data_o[12] )
  );
  NAND _304_ (
    .A(_000_),
    .B(_047_),
    .Y(_133_)
  );
  XOR _305_ (
    .A(_051_),
    .B(_133_),
    .Y(\data_o[13] )
  );
endmodule
